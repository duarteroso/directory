module directory

fn init() {
}
