module vidirectory

fn init() {
}
